module verilog_array_test(
    input [7:0] mem,
    output reg count, 
    output reg [3:0] out
);

    case(mem)
    begin
        8'h00 : count = 4'h0;
        8'h01 : count = 4'h1;
        8'h02 : count = 4'h1;
        8'h03 : count = 4'h2;
        8'h04 : count = 4'h1;
        8'h05 : count = 4'h2;
        8'h06 : count = 4'h2;
        8'h07 : count = 4'h3;
        8'h08 : count = 4'h1;
        8'h09 : count = 4'h1;
        8'h0a : count = 4'h2;
        8'h0b : count = 4'h3;
        8'h0c : count = 4'h2;
        8'h0d : count = 4'h3;
        8'h0e : count = 4'h3;
        8'h0f : count = 4'h4;

        8'h10 : count = 4'h1;
        8'h11 : count = 4'h2;
        8'h12 : count = 4'h2;
        8'h13 : count = 4'h3;
        8'h14 : count = 4'h2;
        8'h15 : count = 4'h3;
        8'h16 : count = 4'h3;
        8'h17 : count = 4'h4;
        8'h18 : count = 4'h2;
        8'h19 : count = 4'h2;
        8'h1a : count = 4'h3;
        8'h1b : count = 4'h4;
        8'h1c : count = 4'h3;
        8'h1d : count = 4'h4;
        8'h1e : count = 4'h4;
        8'h1f : count = 4'h5;

        8'h20 : count = 4'h1;
        8'h21 : count = 4'h2;
        8'h22 : count = 4'h1;
        8'h23 : count = 4'h1;
        8'h24 : count = 4'h1;
        8'h25 : count = 4'h1;
        8'h26 : count = 4'h1;
        8'h27 : count = 4'h1;
        8'h28 : count = 4'h1;
        8'h29 : count = 4'h1;
        8'h2a : count = 4'h1;
        8'h2b : count = 4'h1;
        8'h2c : count = 4'h1;
        8'h2d : count = 4'h1;
        8'h2e : count = 4'h1;
        8'h2f : count = 4'h1;

        8'h30 : count = 4'h0;
        8'h31 : count = 4'h1;
        8'h32 : count = 4'h1;
        8'h33 : count = 4'h1;
        8'h34 : count = 4'h1;
        8'h35 : count = 4'h1;
        8'h36 : count = 4'h1;
        8'h37 : count = 4'h1;
        8'h38 : count = 4'h1;
        8'h39 : count = 4'h1;
        8'h3a : count = 4'h1;
        8'h3b : count = 4'h1;
        8'h3c : count = 4'h1;
        8'h3d : count = 4'h1;
        8'h3e : count = 4'h1;
        8'h3f : count = 4'h1;

        8'h40 : count = 4'h0;
        8'h41 : count = 4'h1;
        8'h42 : count = 4'h1;
        8'h43 : count = 4'h1;
        8'h44 : count = 4'h1;
        8'h45 : count = 4'h1;
        8'h46 : count = 4'h1;
        8'h47 : count = 4'h1;
        8'h48 : count = 4'h1;
        8'h49 : count = 4'h1;
        8'h4a : count = 4'h1;
        8'h4b : count = 4'h1;
        8'h4c : count = 4'h1;
        8'h4d : count = 4'h1;
        8'h4e : count = 4'h1;
        8'h4f : count = 4'h1;

        8'h50 : count = 4'h0;
        8'h51 : count = 4'h1;
        8'h52 : count = 4'h1;
        8'h53 : count = 4'h1;
        8'h54 : count = 4'h1;
        8'h55 : count = 4'h1;
        8'h56 : count = 4'h1;
        8'h57 : count = 4'h1;
        8'h58 : count = 4'h1;
        8'h59 : count = 4'h1;
        8'h5a : count = 4'h1;
        8'h5b : count = 4'h1;
        8'h5c : count = 4'h1;
        8'h5d : count = 4'h1;
        8'h5e : count = 4'h1;
        8'h5f : count = 4'h1;

        8'h60 : count = 4'h0;
        8'h61 : count = 4'h1;
        8'h62 : count = 4'h1;
        8'h63 : count = 4'h1;
        8'h64 : count = 4'h1;
        8'h65 : count = 4'h1;
        8'h66 : count = 4'h1;
        8'h67 : count = 4'h1;
        8'h68 : count = 4'h1;
        8'h69 : count = 4'h1;
        8'h6a : count = 4'h1;
        8'h6b : count = 4'h1;
        8'h6c : count = 4'h1;
        8'h6d : count = 4'h1;
        8'h6e : count = 4'h1;
        8'h6f : count = 4'h1;

        8'h70 : count = 4'h0;
        8'h71 : count = 4'h1;
        8'h72 : count = 4'h1;
        8'h73 : count = 4'h1;
        8'h74 : count = 4'h1;
        8'h75 : count = 4'h1;
        8'h76 : count = 4'h1;
        8'h77 : count = 4'h1;
        8'h78 : count = 4'h1;
        8'h79 : count = 4'h1;
        8'h7a : count = 4'h1;
        8'h7b : count = 4'h1;
        8'h7c : count = 4'h1;
        8'h7d : count = 4'h1;
        8'h7e : count = 4'h1;
        8'h7f : count = 4'h1;

        8'h80 : count = 4'h0;
        8'h81 : count = 4'h1;
        8'h82 : count = 4'h1;
        8'h83 : count = 4'h1;
        8'h84 : count = 4'h1;
        8'h85 : count = 4'h1;
        8'h86 : count = 4'h1;
        8'h87 : count = 4'h1;
        8'h88 : count = 4'h1;
        8'h89 : count = 4'h1;
        8'h8a : count = 4'h1;
        8'h8b : count = 4'h1;
        8'h8c : count = 4'h1;
        8'h8d : count = 4'h1;
        8'h8e : count = 4'h1;
        8'h8f : count = 4'h1;

        8'h90 : count = 4'h0;
        8'h91 : count = 4'h1;
        8'h92 : count = 4'h1;
        8'h93 : count = 4'h1;
        8'h94 : count = 4'h1;
        8'h95 : count = 4'h1;
        8'h96 : count = 4'h1;
        8'h97 : count = 4'h1;
        8'h98 : count = 4'h1;
        8'h99 : count = 4'h1;
        8'h9a : count = 4'h1;
        8'h9b : count = 4'h1;
        8'h9c : count = 4'h1;
        8'h9d : count = 4'h1;
        8'h9e : count = 4'h1;
        8'h9f : count = 4'h1;

        8'ha0 : count = 4'h0;
        8'ha1 : count = 4'h1;
        8'ha2 : count = 4'h1;
        8'ha3 : count = 4'h1;
        8'ha4 : count = 4'h1;
        8'ha5 : count = 4'h1;
        8'ha6 : count = 4'h1;
        8'ha7 : count = 4'h1;
        8'ha8 : count = 4'h1;
        8'ha9 : count = 4'h1;
        8'haa : count = 4'h1;
        8'hab : count = 4'h1;
        8'hac : count = 4'h1;
        8'had : count = 4'h1;
        8'hae : count = 4'h1;
        8'haf : count = 4'h1;

        8'hb0 : count = 4'h0;
        8'hb1 : count = 4'h1;
        8'hb2 : count = 4'h1;
        8'hb3 : count = 4'h1;
        8'hb4 : count = 4'h1;
        8'hb5 : count = 4'h1;
        8'hb6 : count = 4'h1;
        8'hb7 : count = 4'h1;
        8'hb8 : count = 4'h1;
        8'hb9 : count = 4'h1;
        8'hba : count = 4'h1;
        8'hbb : count = 4'h1;
        8'hbc : count = 4'h1;
        8'hbd : count = 4'h1;
        8'hbe : count = 4'h1;
        8'hbf : count = 4'h1;

        8'hc0 : count = 4'h0;
        8'hc1 : count = 4'h1;
        8'hc2 : count = 4'h1;
        8'hc3 : count = 4'h1;
        8'hc4 : count = 4'h1;
        8'hc5 : count = 4'h1;
        8'hc6 : count = 4'h1;
        8'hc7 : count = 4'h1;
        8'hc8 : count = 4'h1;
        8'hc9 : count = 4'h1;
        8'hca : count = 4'h1;
        8'hcb : count = 4'h1;
        8'hcc : count = 4'h1;
        8'hcd : count = 4'h1;
        8'hce : count = 4'h1;
        8'hcf : count = 4'h1;

        8'hh0 : count = 4'h0;
        8'hh1 : count = 4'h1;
        8'hh2 : count = 4'h1;
        8'hh3 : count = 4'h1;
        8'hh4 : count = 4'h1;
        8'hh5 : count = 4'h1;
        8'hh6 : count = 4'h1;
        8'hh7 : count = 4'h1;
        8'hh8 : count = 4'h1;
        8'hh9 : count = 4'h1;
        8'hha : count = 4'h1;
        8'hhb : count = 4'h1;
        8'hhc : count = 4'h1;
        8'hhd : count = 4'h1;
        8'hhe : count = 4'h1;
        8'hhf : count = 4'h1;

        8'he0 : count = 4'h0;
        8'he1 : count = 4'h1;
        8'he2 : count = 4'h1;
        8'he3 : count = 4'h1;
        8'he4 : count = 4'h1;
        8'he5 : count = 4'h1;
        8'he6 : count = 4'h1;
        8'he7 : count = 4'h1;
        8'he8 : count = 4'h1;
        8'he9 : count = 4'h1;
        8'hea : count = 4'h1;
        8'heb : count = 4'h1;
        8'hec : count = 4'h1;
        8'hed : count = 4'h1;
        8'hee : count = 4'h1;
        8'hef : count = 4'h1;

        8'hf0 : count = 4'h0;
        8'hf1 : count = 4'h1;
        8'hf2 : count = 4'h1;
        8'hf3 : count = 4'h1;
        8'hf4 : count = 4'h1;
        8'hf5 : count = 4'h1;
        8'hf6 : count = 4'h1;
        8'hf7 : count = 4'h1;
        8'hf8 : count = 4'h1;
        8'hf9 : count = 4'h1;
        8'hfa : count = 4'h1;
        8'hfb : count = 4'h1;
        8'hfc : count = 4'h1;
        8'hfd : count = 4'h1;
        8'hfe : count = 4'h1;
        8'h0f : count = 4'h1;

        default : count = 4'h0;
    endcase
endmodule