module shift_right_8(
    input [7:0] ip,
    input load,
    input shift,
    input clk,
    input clr,
    output reg shift_out,
);

